/***********************************************************************
 * A SystemVerilog testbench for an instruction register; This file
 * contains the interface to connect the testbench to the design
 **********************************************************************/
interface tb_ifc (input logic clk);
  timeunit 1ns/1ns;

  // user-defined types are defined in instr_register_pkg.sv
  import instr_register_pkg::*;

  // ADD CODE TO DECLARE THE INTERFACE SIGNALS

modport dut (input load_en, reset_n, operand_a,operand_b, opcode, write_pointer,read_pointer
            output instruction_word);

modport test (input load_en, reset_n, operand_a,operand_b, opcode, write_pointer,read_pointer
            output instruction_word);
  
endinterface: tb_ifc

